`include "adder.v" 
`include "alu.v"
`include "d_ff.v" 
`include "control_unit.v" 
`include "counter.v" 
`include "full-adder.v" 
`include "mod4-count.v"
`include "mux2-1-8bit.v" 
`include "mux2-1.v" 
`include "complement.v"
`include "mux4-1.v"
`include "mux4-1-8bit.v" 
`include "shift_reg_lr.v"
`include "sr_ff.v"