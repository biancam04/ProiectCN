// Booth Multiplier Structural Datapath (Fixed)
module booth_datapath (
    input wire clk,
    input wire reset,
    input wire start,
    input wire [7:0] multiplicand,  // inbus_b
    input wire [7:0] multiplier,    // inbus_a
    output reg [15:0] product,
    output wire done
);
    reg [7:0] A, M, Q;
    reg Q_1;
    reg [3:0] count;
    reg busy;

    // Assign done signal
    assign done = ~busy;

    // State machine logic
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            A <= 8'b0;
            Q <= 8'b0;
            M <= 8'b0;
            Q_1 <= 1'b0;
            count <= 4'd0;
            busy <= 1'b0;
            product <= 16'b0;
        end else begin
            if (start) begin
                A <= 8'b0;
                Q <= multiplier;
                M <= multiplicand;
                Q_1 <= 1'b0;
                count <= 4'd8;
                busy <= 1'b1;
                product <= 16'b0;
            end else if (busy) begin
                case ({Q[0], Q_1})
                    2'b01: A <= A + M;  // A = A + M
                    2'b10: A <= A - M;  // A = A - M
                    default: A <= A;    // No operation
                endcase

                // Arithmetic right shift {A, Q, Q-1}
                {A, Q, Q_1} <= {A[7], A, Q};

                count <= count - 1;
                if (count == 4'd1) begin
                    busy <= 1'b0;  // Finished after 8 shifts
                    product <= {A, Q};
                end
            end
        end
    end

endmodule

