library verilog;
use verilog.vl_types.all;
entity alu_top_tb is
end alu_top_tb;
