module counter (
    input  wire clk,     // Clock input
    input  wire rst,     // Active-high synchronous reset
    input  wire en,      // Enable counting
    output reg  [2:0] o  // 3-bit count output
);

    always @(posedge clk) begin
        if (rst)
            o <= 3'b000;
        else if (en)
            o <= o + 1;
    end

endmodule
